`include "uvm_hdrs.sv"
`include "eth_pkt.sv"
`include "top.sv"
