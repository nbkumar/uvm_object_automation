import uvm_pkg::*;
`include "uvm_macros.svh"
